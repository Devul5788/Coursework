/*

	Module: finalProject.sv
	Authors: Shubham & Devul

*/

module finalProject (

      ///////// Clocks /////////
      input     MAX10_CLK1_50, 

      ///////// KEY /////////
      input    [ 1: 0]   KEY,

      ///////// SW /////////
      input    [ 9: 0]   SW,

      ///////// LEDR /////////
      output   [ 9: 0]   LEDR,

      ///////// HEX /////////
      output   [ 7: 0]   HEX0,
      output   [ 7: 0]   HEX1,
      output   [ 7: 0]   HEX2,
      output   [ 7: 0]   HEX3,
      output   [ 7: 0]   HEX4,
      output   [ 7: 0]   HEX5,

      ///////// SDRAM /////////
      output             DRAM_CLK,
      output             DRAM_CKE,
      output   [12: 0]   DRAM_ADDR,
      output   [ 1: 0]   DRAM_BA,
      inout    [15: 0]   DRAM_DQ,
      output             DRAM_LDQM,
      output             DRAM_UDQM,
      output             DRAM_CS_N,
      output             DRAM_WE_N,
      output             DRAM_CAS_N,
      output             DRAM_RAS_N,

      ///////// VGA /////////
      output             VGA_HS,
      output             VGA_VS,
      output   [ 3: 0]   VGA_R,
      output   [ 3: 0]   VGA_G,
      output   [ 3: 0]   VGA_B,


      ///////// ARDUINO /////////
      inout    [15: 0]   ARDUINO_IO,
      inout              ARDUINO_RESET_N, 

		input [18:0] addressFromPi,
		output dataToPi, restartToPi, charDoneToPi, solveToPi,
		input answerReadyFromPi
);


// Local variables

logic [18:0] answer;

always_comb begin
	answer = 0;
	if(answerReadyFromPi == 1) begin
		answer = addressFromPi;
	end
end

logic Reset_h, vssig, blank, sync, VGA_Clk;


//=======================================================
//  REG/WIRE declarations
//=======================================================
	logic SPI0_CS_N, SPI0_SCLK, SPI0_MISO, SPI0_MOSI, USB_GPX, USB_IRQ, USB_RST;
	logic [3:0] hex_num_4, hex_num_3, hex_num_1, hex_num_0; //4 bit input hex digits
	logic [1:0] signs;
	logic [1:0] hundreds;
	logic [9:0] drawxsig, drawysig, ballxsig, ballysig, ballsizesig;
	logic [7:0] Red, Blue, Green;
	logic [7:0] keycode;
	logic [7:0] mousebutton;
	logic [31:0] mousex;
	logic [31:0] mousey;

//=======================================================
//  Structural coding
//=======================================================
	assign ARDUINO_IO[10] = SPI0_CS_N;
	assign ARDUINO_IO[13] = SPI0_SCLK;
	assign ARDUINO_IO[11] = SPI0_MOSI;
	assign ARDUINO_IO[12] = 1'bZ;
	assign SPI0_MISO = ARDUINO_IO[12];
	
	assign ARDUINO_IO[9] = 1'bZ; 
	assign USB_IRQ = ARDUINO_IO[9];
		
	//Assignments specific to Circuits At Home UHS_20
	assign ARDUINO_RESET_N = USB_RST;
	assign ARDUINO_IO[7] = USB_RST;//USB reset 
	assign ARDUINO_IO[8] = 1'bZ; //this is GPX (set to input)
	assign USB_GPX = 1'b0;//GPX is not needed for standard USB host - set to 0 to prevent interrupt
	
	//Assign uSD CS to '1' to prevent uSD card from interfering with USB Host (if uSD card is plugged in)
	assign ARDUINO_IO[6] = 1'b1;
	
	//HEX drivers to convert numbers to HEX output
	
	//	HexDriver hex_driver0 (addressFromPi[3:0], HEX0[6:0]);
	//	HexDriver hex_driver1 (addressFromPi[7:4], HEX1[6:0]);
	//	HexDriver hex_driver2 (addressFromPi[11:8], HEX2[6:0]);
	//	HexDriver hex_driver3 (addressFromPi[15:12], HEX3[6:0]);
	//	HexDriver hex_driver4 (addressFromPi[18:16], HEX4[6:0]);

	HexDriver hex_driver0 (answer[3:0], HEX0[7:0]);
	HexDriver hex_driver1 (answer[7:4], HEX1[7:0]);
	HexDriver hex_driver2 (answer[11:8], HEX2[7:0]);
	SignDriver hex_driver3 (answer[18], HEX3[7:0]);
	
	HexDriver hex_driver4 (addressFromPi[15:12], HEX4[7:0]);
	HexDriver hex_driver5 (addressFromPi[18:16], HEX5[7:0]);
	
	//Assign one button to reset
	assign {Reset_h}=~ (KEY[0]);

	//Our A/D converter is only 12 bit
	assign VGA_R = Red[7:4];
	assign VGA_B = Blue[7:4];
	assign VGA_G = Green[7:4];
	
	
	final_project_soc u0(
		.clk_clk                           (MAX10_CLK1_50),  //clk.clk
		.reset_reset_n                     (1'b1),           //reset.reset_n
		.altpll_0_locked_conduit_export    (),               //altpll_0_locked_conduit.export
		.altpll_0_phasedone_conduit_export (),               //altpll_0_phasedone_conduit.export
		.altpll_0_areset_conduit_export    (),               //altpll_0_areset_conduit.export
		.key_external_connection_export    (KEY),            //key_external_connection.export

		//SDRAM
		.sdram_clk_clk(DRAM_CLK),                            //clk_sdram.clk
		.sdram_wire_addr(DRAM_ADDR),                         //sdram_wire.addr
		.sdram_wire_ba(DRAM_BA),                             //.ba
		.sdram_wire_cas_n(DRAM_CAS_N),                       //.cas_n
		.sdram_wire_cke(DRAM_CKE),                           //.cke
		.sdram_wire_cs_n(DRAM_CS_N),                         //.cs_n
		.sdram_wire_dq(DRAM_DQ),                             //.dq
		.sdram_wire_dqm({DRAM_UDQM,DRAM_LDQM}),              //.dqm
		.sdram_wire_ras_n(DRAM_RAS_N),                       //.ras_n
		.sdram_wire_we_n(DRAM_WE_N),                         //.we_n

		//USB SPI	
		.spi0_SS_n(SPI0_CS_N),
		.spi0_MOSI(SPI0_MOSI),
		.spi0_MISO(SPI0_MISO),
		.spi0_SCLK(SPI0_SCLK),
		
		//USB GPIO
		.usb_rst_export(USB_RST),
		.usb_irq_export(USB_IRQ),
		.usb_gpx_export(USB_GPX),
		
		//LEDs and HEX
		.keycode_export(keycode),
		.mousebutton_export(mousebutton),
		.mousex_export(mousex),
		.mousey_export(mousey)
	 );


	vga_controller myVGA (.Clk(MAX10_CLK1_50),    
								 .Reset(Reset_h),     	 
								 .hs(VGA_HS),        	 
								 .vs(VGA_VS),        	 
								 .pixel_clk(VGA_Clk), 	 
								 .blank(blank),     		 
								 .sync(sync),     		 
								 .DrawX(drawxsig),     	 
								 .DrawY(drawysig));   	 

	
	cursor myCursor(.Reset(Reset_h), 
						 .frame_clk(VGA_VS),
						 .keycode(keycode),
						 .BallX(ballxsig), 
						 .BallY(ballysig), 
						 .BallS(ballsizesig),
						 .mouseX(mousex),
						 .mouseY(mousey),
						 .mouseButton(mousebutton));
	
	canvas myCanvas(.BallX(ballxsig), 
						 .BallY(ballysig),
						 .mouseButton(mousebutton), 
						 .DrawX(drawxsig), 
						 .DrawY(drawysig), 
						 .Ball_size(ballsizesig),
						 .Red(Red), 
						 .Green(Green),
						 .Blue(Blue),
						 .blank(blank),
						 .pixel_clk(VGA_Clk),
						 .clk(MAX10_CLK1_50),
						 .addressFromPi(addressFromPi),
						 .dataToPi(dataToPi),
						 .restartToPi(restartToPi),
						 .charDoneToPi(charDoneToPi),
						 .solveToPi(solveToPi),
						 .LEDR(LEDR),
						 .SW(SW),
						 .answerReadyFromPi(answerReadyFromPi));

endmodule
