/* MODIFY. Your cache design. It contains the cache
controller, cache datapath, and bus adapter. */

module cache #(
    parameter s_offset = 5,
    parameter s_index  = 3,
    parameter s_tag    = 32 - s_offset - s_index,
    parameter s_mask   = 2**s_offset,
    parameter s_line   = 8*s_mask,
    parameter num_sets = 2**s_index
)
(
    input clk,
    input rst,

    /* CPU memory signals */
    input   logic [31:0]    mem_address,        //The memory system is accessed using this 32 bit signal. 
                                                //It specifies the address that is to be read or written.
    output  logic [31:0]    mem_rdata,          //32-bit data bus for receiving data from the memory system.
    input   logic [31:0]    mem_wdata,          //32-bit data bus for sending data to the memory system.
    input   logic           mem_read,           //Active high signal that tells the memory system that the 
                                                //address is valid and the processor is trying to perform a memory read.
    input   logic           mem_write,          //Active high signal that tells the memory system that the address is 
                                                //valid and the processor is trying to perform a memory write.
    input   logic [3:0]     mem_byte_enable,    //A mask describing which byte(s) of memory should be written on a memory write. 
                                                //4'b0000 -> Don't write to memory even if write_enable is 1. 
                                                //4'b???? -> Write only bytes specified if the bit is 1.
                                                //4'b1111 -> Write all bytes of a word to memory when mem_write becomes active
    output  logic           mem_resp,           //Active high signal generated by the memory system indicating that the memory has
                                                //finished the requested operation.

    /* Physical memory signals */
    output  logic [31:0]    pmem_address,       //Physical memory is accessed using this 32-bit signal. It specifies the physical 
                                                //memory address that is to be read or written.
    input   logic [255:0]   pmem_rdata,         //256-bit data bus for receiving data from physical memory.
    output  logic [255:0]   pmem_wdata,         //256-bit data bus for sending data to physical memory.
    output  logic           pmem_read,          //Active high signal that tells the memory interface that the address 
                                                //is valid and the cache is trying to perform a physical memory read.
    output  logic           pmem_write,         //Active high signal that tells the memory interface that the address
                                                //is valid and the cache is trying to perform a physical memory write.
    input   logic           pmem_resp           //Active high signal generated by the memory interface indicating
                                                //that the memory operation has completed.
);

// load signals for arrays
logic dirty_load0;
logic dirty_load1;
logic valid_load0;
logic valid_load1;
logic lru_load;
logic tag_load0;
logic tag_load1;

// input signals for arrays
logic lru_input;
logic dirty_input0;
logic dirty_input1;
logic valid_input0;
logic valid_input1;

// output signals for arrays
logic dirty_out0;
logic dirty_out1;
logic valid_out0;
logic valid_out1;
logic lru_out;

// set associative signals
logic hit0;
logic hit1;
logic way_select0;
logic way_select1;

// internal signals for datapath
logic [255:0] mem_wdata256; 
logic [31:0] mem_byte_enable256; 
logic [255:0] mem_rdata256; 
logic [31:0] address;
logic pmem_addr_sel;
assign address = mem_address;

// signals for data byte enable when writing
logic [31:0] mem_byte_enable256_0;
logic [31:0] mem_byte_enable256_1;

cache_control control
(.*);

cache_datapath datapath
(.*);

bus_adapter bus_adapter
(.*);

endmodule : cache
